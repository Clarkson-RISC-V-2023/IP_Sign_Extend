module <new_ip_name> # (
    // Parameters go here
)(
    // Define ports, inputs and outputs
);

    // Define regs & wires

    // Define RTL

endmodule